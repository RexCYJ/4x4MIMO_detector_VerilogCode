`timescale 1ns / 1ps

`include "parameters.v"

module InnerProduct(

    );
    
    
    
endmodule
